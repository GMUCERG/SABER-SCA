--------------------------------------------------------------------------------
--! @file       decaps_tv_shared_pkg_2.vhd
--! @author     Abubakr Abdulgadir
--! @copyright  Copyright (c) 2021 Cryptographic Engineering Research Group
--!             ECE Department, George Mason University Fairfax, VA, U.S.A.
--!             All rights Reserved.
--------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.all;
use ieee.numeric_std.all;

use work.saber_pkg.all;
use work.saber_pr_pkg.all;

package decaps_tv_shared_pkg_2 is


    type decaps_input_shared_arr_type is array (0 to 2**DIN_FIFO_LOG2DEPTH-1) of std_logic_vector(DIN_FIFO_WIDTH-1 downto 0);
    constant DECAPS_INPUT_DATA : decaps_input_shared_arr_type := 
    (
    --opcode =================================================================================================
    OPCODE_DECAPS,
    --PK======================================================================================================
    --b polycev
    x"aa45", x"77e7", x"b8f8", x"aa90", x"0420", x"9891", x"b38d", x"e401", x"0b78", x"58eb", x"1278", x"98cd", x"9f14", x"3363", x"02dd", x"75b9", x"4f99", x"d675", x"afc8", x"2986", x"0061", x"6bd3", x"483e", x"30ff", x"93ff", x"27d7", x"9126", x"9253", x"7e9d", x"795d", x"962a", x"d662", x"e046", x"05ef", x"f8ef", x"e65c", x"3df5", x"f833", x"7668", x"f2e7", x"f274", x"6e04", x"12f2", x"03c1", x"3f96", x"4bba", x"eaf6", x"1c77", x"af40", x"e173", x"735c", x"98cb", x"3158", x"b0f2", x"b8d8", x"4f5f", x"1990", x"835c", x"7c6d", x"d411", x"98c0", x"5a56", x"af01", x"70cf", x"2b17", x"a4af", x"a47d", x"e427", x"7434", x"9346", x"b4ff", x"a54d", x"721c", x"9e6c", x"6600", x"944f", x"e380", x"a776", x"c7ca", x"22a2", x"488b", x"82b6", x"6fd2", x"e50a", x"8672", x"5d9c", x"f5f2", x"602b", x"1585", x"3968", x"c1c7", x"583a", x"9775", x"8798", x"41b0", x"bda4", x"6976", x"0e35", x"92f7", x"163c", x"a5c5", x"c83a", x"4fe3", x"84af", x"d123", x"672e", x"f23a", x"30bd", x"6413", x"989d", x"8a68", x"60eb", x"bf89", x"8a3a", x"a505", x"6f8a", x"5cb9", x"8b04", x"4aac", x"78a7", x"ab0f", x"5486", x"5a0c", x"79a2", x"f943", x"e9d9", x"1ff7", x"fa2c", x"d2f0", x"8d61", x"688e", x"8de2", x"eb33", x"23d8", x"c791", x"7e92", x"24d7", x"06cc", x"a540", x"3d6b", x"ee3e", x"9b81", x"52fa", x"0ed0", x"a347", x"801d", x"c6c4", x"9ea6", x"3fd9", x"f747", x"9f73", x"bd6e", x"6216", x"5013", x"8233", x"6aef", x"c2da", x"1f91", x"2b9a", x"0cf0", x"837f", x"1cce", x"933e", x"a910", x"602b", x"a3f8", x"1d03", x"ed2d", x"5e1d", x"ff59", x"04dc", x"66cd", x"3cd1", x"c29e", x"3949", x"f35d", x"096c", x"db48", x"d785", x"4327", x"955c", x"e9b7", x"b7fe", x"d11e", x"97b7", x"26fb", x"d519", x"324f", x"6947", x"797b", x"a27e", x"d26d", x"3a17", x"d9de", x"0cdf", x"f7a4", x"7e75", x"80fb", x"07ac", x"b053", x"0651", x"eabe", x"54e6", x"9001", x"f3a9", x"9907", x"55fe", x"94a0", x"faa5", x"4545", x"7d7a", x"36b0", x"ced8", x"21f3", x"1d58", x"ef7e", x"d8fc", x"8e72", x"42d8", x"4eec", x"d69f", x"5f41", x"35c4", x"e893", x"6e2f", x"7b1d", x"53e4", x"f424", x"d007", x"7cd0", x"7668", x"e77d", x"db30", x"0e0c", x"bf8f", x"c65c", x"161e", x"6e28", x"f76d", x"1ed6", x"001a", x"2f76", x"ae0c", x"cf41", x"17bb", x"9080", x"5e9d", x"bdc2", x"31bb", x"0eab", x"fdae", x"16a9", x"6339", x"cd46", x"e3a3", x"77e5", x"f1e3", x"60a1", x"8bad", x"8c69", x"37bd", x"01b7", x"5e2a", x"c383", x"38fb", x"5073", x"5492", x"a7bb", x"65a0", x"9e9c", x"4521", x"5489", x"98f9", x"4c28", x"34df", x"c235", x"e75f", x"58a0", x"52c2", x"bf53", x"4342", x"786e", x"1141", x"c693", x"82be", x"0c8e", x"9316", x"946b", x"9a28", x"7716", x"0e76", x"125f", x"824e", x"50a5", x"ed47", x"14e1", x"22a1", x"8e49", x"91e6", x"9899", x"7cc6", x"284d", x"5c3b", x"6d17", x"2339", x"9649", x"9e6f", x"0030", x"29c5", x"4bf5", x"9b43", x"0474", x"f282", x"bddd", x"7d80", x"cb61", x"3642", x"afab", x"3b88", x"7b0a", x"c5ad", x"c208", x"384d", x"f8b1", x"dba0", x"307c", x"8247", x"0fce", x"1f40", x"5011", x"babc", x"8fe8", x"2f57", x"e71d", x"9eb5", x"d1c5", x"3fb7", x"defb", x"1f26", x"3315", x"b76a", x"1765", x"f24d", x"aab4", x"c7cf", x"e506", x"02c7", x"9f59", x"5197", x"1798", x"2679", x"d8f7", x"f5c1", x"56b0", x"cd4a", x"4553", x"4277", x"524e", x"adbc", x"22b7", x"22c0", x"5a4c", x"b571", x"4f09", x"1ac1", x"9636", x"7e30", x"ae05", x"9ae6", x"8b93", x"6c52", x"7a29", x"ef3d", x"cc41", x"39e3", x"fa00", x"ea52", x"3fa6", x"a2a0", x"e2b5", x"47d5", x"1017", x"21c4", x"6647", x"b747", x"5c83", x"005c", x"f04a", x"e5c7", x"f10e", x"3686", x"5e69", x"d834", x"0569", x"129a", x"ee96", x"50ea", x"0c79", x"537a", x"a5df", x"1cfd", x"d252", x"c6f0", x"d8b3", x"f8b8", x"b11d", x"f561", x"7431", x"f134", x"e31f", x"a67b", x"7dba", x"fff3", x"7ab7", x"c1f5", x"7f32", x"35c4", x"9131", x"020d", x"f48b", x"98fe", x"b189", x"c562", x"7225", x"acec", x"8d05", x"93b3", x"d9f3", x"79d8", x"36b4", x"1425", x"1ade", x"452a", x"0ca2", x"ffff", x"592c", x"82d4", x"a8e0", x"5e45", x"b7a4", x"97e7", x"f1eb", x"ae50", x"c854", x"4aa1", x"6ae1", x"b045", x"2fa9", x"b8e5", x"a5d9", x"7124", x"b54e", x"9cf6", x"87c5", x"134c", x"7619", x"ed02", x"f555", x"3135", x"7305", x"5a95", x"30d0", x"fae5", x"77df", x"f4e1", x"4058", x"d488", x"c7ad", x"a4eb", x"6984", x"a07a", x"4e5b", x"a618", x"0335", x"8f11", x"6467", x"75e2", x"fc7e", x"2880", x"91fc", 
    --SEED_A
    x"6236", x"0808", x"1330", x"04de", x"4a63", x"8f4e", x"2bfd", x"6486", x"d98c", x"cd8e", x"c674", x"26f4", x"af2d", x"622f", x"bc8b", x"c48b",
    --SEED_A second share (no need to share but this is just a work around since SHA3 needs 2 shares).
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000",
    --END_PK===================================================================================================
    
    --SK--share0=======================================================================================================
    --S polyvec 
       --orig
--    x"0001",x"1fff",x"0000",x"0000",x"1ffe",x"0002",x"0001",x"0000",x"1fff",x"0001",x"0000",x"0001",x"1ffe",x"1fff",x"0003",x"1fff",x"1ffe",x"1ffd",x"1fff",x"0003",x"0001",x"0002",x"0000",x"0001",x"0002",x"0002",x"1fff",x"0000",x"0000",x"1fff",x"0001",x"0000",x"1ffe",x"0000",x"1ffc",x"0000",x"0001",x"0000",x"1fff",x"0000",x"1fff",x"0001",x"0000",x"1ffe",x"1ffd",x"0000",x"1ffe",x"1ffd",x"1fff",x"1fff",x"1fff",x"0000",x"1fff",x"1fff",x"1ffe",x"0001",x"0000",x"0000",x"1fff",x"1fff",x"0000",x"0001",x"0001",x"0002",x"0000",x"0001",x"0001",x"0002",x"1fff",x"0000",x"0000",x"0000",x"0001",x"0001",x"0001",x"0003",x"0001",x"0001",x"1fff",x"1fff",x"1ffd",x"0001",x"1fff",x"0001",x"1fff",x"0000",x"1ffe",x"0001",x"1fff",x"0001",x"1ffe",x"0000",x"1ffe",x"1ffe",x"0001",x"0000",x"0000",x"0000",x"0000",x"0001",x"0001",x"1fff",x"1fff",x"0000",x"0001",x"0000",x"1fff",x"0001",x"0001",x"1ffd",x"1ffe",x"0000",x"0003",x"1ffe",x"0000",x"0002",x"1ffe",x"0000",x"0001",x"0003",x"0000",x"0001",x"0001",x"0001",x"1fff",x"1ffd",x"1ffe",x"0000",x"1ffe",x"0000",x"0001",x"1fff",x"1fff",x"1ffe",x"0001",x"0000",x"1fff",x"0002",x"1fff",x"0000",x"0004",x"0001",x"1ffe",x"0003",x"1fff",x"0002",x"0001",x"0002",x"0003",x"0000",x"1fff",x"0000",x"0000",x"1ffe",x"1fff",x"0000",x"1fff",x"0000",x"0002",x"1fff",x"0001",x"0001",x"1ffe",x"1fff",x"1ffd",x"0000",x"0002",x"0000",x"0002",x"0000",x"0002",x"0001",x"1ffe",x"1fff",x"1ffe",x"0000",x"0000",x"1fff",x"0003",x"1ffe",x"0000",x"0000",x"1ffe",x"0001",x"0001",x"0001",x"0001",x"0000",x"0000",x"0000",x"0002",x"1fff",x"1fff",x"0001",x"0000",x"0001",x"1fff",x"0001",x"0000",x"0001",x"1ffd",x"1ffe",x"0000",x"0000",x"1ffe",x"1fff",x"1fff",x"0000",x"0001",x"0001",x"1fff",x"0001",x"0001",x"0002",x"1ffe",x"1ffe",x"0001",x"1ffe",x"0002",x"0000",x"1ffe",x"0001",x"1fff",x"0000",x"1fff",x"1fff",x"0001",x"1fff",x"1ffe",x"0002",x"1ffe",x"0001",x"0001",x"0000",x"0000",x"1fff",x"0000",x"1fff",x"1fff",x"0001",x"0002",x"0001",x"1fff",x"0000",x"0001",x"0002",x"1fff",x"0001",x"0002",x"0001",x"0001",x"1fff",x"0000",x"0000",x"1fff",x"0001",
--    x"1fff",x"0000",x"0000",x"0001",x"1fff",x"0000",x"0000",x"0001",x"0003",x"1fff",x"0001",x"0000",x"0001",x"0000",x"1ffe",x"0001",x"0001",x"0001",x"1ffe",x"1fff",x"0002",x"1fff",x"1ffd",x"0001",x"1fff",x"0001",x"0000",x"0000",x"0001",x"0003",x"1ffe",x"1ffd",x"0000",x"0000",x"0000",x"1fff",x"0000",x"1ffe",x"0000",x"0001",x"0000",x"0000",x"0000",x"0000",x"0001",x"0002",x"0000",x"0001",x"1ffd",x"0000",x"1fff",x"0002",x"1ffe",x"1ffe",x"0002",x"0001",x"0001",x"0002",x"0002",x"0000",x"1ffe",x"0000",x"0000",x"1ffe",x"0001",x"0001",x"0001",x"0002",x"0001",x"0001",x"0001",x"1ffe",x"0000",x"0001",x"0002",x"1fff",x"0002",x"0002",x"1fff",x"1fff",x"1fff",x"0003",x"0000",x"0000",x"1ffe",x"0001",x"0000",x"0000",x"0000",x"0001",x"0000",x"0001",x"0000",x"1fff",x"1fff",x"0000",x"0001",x"0001",x"1fff",x"1fff",x"0000",x"1ffe",x"0002",x"1fff",x"1ffe",x"0000",x"1fff",x"0002",x"0002",x"0000",x"0000",x"0000",x"0000",x"0000",x"1fff",x"0000",x"0000",x"0001",x"0000",x"1fff",x"0000",x"0000",x"0002",x"0001",x"0001",x"1fff",x"0001",x"0001",x"0000",x"0003",x"1fff",x"0001",x"0003",x"1fff",x"1fff",x"0002",x"0000",x"0000",x"0001",x"0000",x"1fff",x"0003",x"0000",x"1ffe",x"1ffe",x"0000",x"1ffe",x"0002",x"0001",x"1ffd",x"0002",x"0001",x"0001",x"1fff",x"0000",x"0000",x"0000",x"1fff",x"0001",x"0001",x"1ffe",x"0002",x"0002",x"1fff",x"0003",x"0001",x"0000",x"0000",x"0002",x"0001",x"0001",x"1ffe",x"1fff",x"0001",x"0001",x"0000",x"0000",x"1fff",x"0001",x"1fff",x"1ffd",x"0002",x"1fff",x"1ffe",x"1fff",x"1ffe",x"0001",x"1ffd",x"0001",x"0001",x"0002",x"0000",x"0001",x"0001",x"0000",x"0000",x"0001",x"1fff",x"1fff",x"1fff",x"0001",x"0001",x"0000",x"0003",x"0001",x"0000",x"0000",x"0000",x"1fff",x"0000",x"0002",x"1fff",x"1ffe",x"0001",x"1fff",x"0002",x"0000",x"0002",x"0002",x"0001",x"0001",x"1ffd",x"0000",x"0001",x"0000",x"0000",x"0000",x"0002",x"0000",x"0001",x"0001",x"0002",x"0000",x"0000",x"0001",x"0001",x"0000",x"1fff",x"1fff",x"0001",x"0000",x"0002",x"1ffe",x"0004",x"1fff",x"1ffe",x"1fff",x"1ffe",x"0000",x"1fff",x"0002",x"0001",x"0001",x"1fff",x"0000",x"1ffe",
--    x"1ffe",x"0000",x"0002",x"1fff",x"0000",x"1ffe",x"1ffe",x"1ffe",x"0000",x"0002",x"0000",x"1fff",x"1fff",x"1fff",x"0001",x"0000",x"0002",x"0003",x"0000",x"1ffe",x"0001",x"1ffd",x"0002",x"0002",x"0001",x"0001",x"1fff",x"1fff",x"1fff",x"0000",x"0000",x"0000",x"0000",x"0000",x"0001",x"0001",x"0001",x"1ffe",x"1ffe",x"1fff",x"0000",x"0002",x"1ffd",x"0001",x"0000",x"0001",x"0001",x"0001",x"1fff",x"1fff",x"0001",x"1ffd",x"0002",x"1fff",x"1fff",x"1ffe",x"1fff",x"0002",x"0000",x"1ffe",x"0001",x"0001",x"1fff",x"0001",x"1ffc",x"1fff",x"0001",x"0002",x"0001",x"0000",x"0000",x"1fff",x"0001",x"0000",x"0001",x"0000",x"1ffe",x"0001",x"1ffd",x"0001",x"0001",x"0000",x"1fff",x"1ffe",x"0001",x"1fff",x"0002",x"1fff",x"1ffe",x"0000",x"0002",x"1ffe",x"0000",x"1fff",x"0000",x"0001",x"0001",x"1ffc",x"0002",x"1fff",x"1ffe",x"0001",x"0001",x"0001",x"0001",x"0000",x"1fff",x"1fff",x"0000",x"1fff",x"1ffe",x"0000",x"1ffe",x"0001",x"0003",x"0000",x"1ffe",x"0002",x"0000",x"1fff",x"0000",x"1fff",x"0000",x"1fff",x"1ffe",x"0002",x"1ffe",x"1fff",x"1fff",x"0002",x"1ffe",x"0000",x"1ffd",x"1fff",x"0000",x"1ffd",x"0001",x"0001",x"1fff",x"1fff",x"0000",x"0000",x"1fff",x"1ffe",x"1ffe",x"0001",x"1ffd",x"0001",x"1ffe",x"1ffe",x"1fff",x"1fff",x"0001",x"1fff",x"0000",x"0001",x"0000",x"0000",x"0000",x"1fff",x"0000",x"0001",x"0002",x"0001",x"1fff",x"0003",x"0001",x"0001",x"0001",x"0001",x"1ffe",x"0000",x"1ffe",x"1fff",x"0000",x"1ffe",x"1ffe",x"1fff",x"1fff",x"1fff",x"0001",x"0000",x"0001",x"1fff",x"0001",x"0001",x"0001",x"0000",x"1fff",x"0000",x"0001",x"0001",x"1fff",x"0001",x"1fff",x"0002",x"0001",x"0002",x"0000",x"0001",x"1ffe",x"0001",x"0001",x"0000",x"0001",x"0001",x"0000",x"1ffe",x"0002",x"0001",x"0000",x"0002",x"0003",x"1fff",x"0001",x"0000",x"0000",x"0001",x"0001",x"0001",x"0001",x"0000",x"0002",x"0000",x"1fff",x"0001",x"1ffe",x"0002",x"0001",x"1fff",x"0000",x"0001",x"0000",x"1ffe",x"1fff",x"1fff",x"1ffe",x"1ffe",x"1fff",x"1ffe",x"0002",x"0000",x"1fff",x"1ffe",x"0000",x"1ffe",x"1fff",x"0001",x"1fff",x"1fff",x"0001",x"0000",x"1fff",x"1ffe",x"0001",x"0002",
    --rand shared
    x"0001",x"0001",x"1fff",x"0000",x"0002",x"0000",x"0000",x"1fff",x"1ffe",x"1fff",x"1fff",x"1fff",x"0000",x"1fff",x"0003",x"0001",x"0000",x"0001",x"0002",x"0001",x"0000",x"0000",x"0000",x"0000",x"1ffe",x"0001",x"1ffd",x"0001",x"1fff",x"0000",x"0002",x"0000",x"1ffe",x"1ffe",x"0000",x"0001",x"0000",x"0000",x"0002",x"0001",x"1ffe",x"1ffe",x"1fff",x"1fff",x"0002",x"1fff",x"1fff",x"1ffd",x"0003",x"0000",x"1fff",x"0002",x"0001",x"1ffe",x"0000",x"1fff",x"0000",x"0001",x"0000",x"1fff",x"0002",x"1ffe",x"0001",x"1ffe",x"1fff",x"0002",x"1ffe",x"0002",x"1ffd",x"0002",x"0000",x"0001",x"1fff",x"0000",x"0002",x"0002",x"1fff",x"0000",x"0001",x"0002",x"1fff",x"1ffe",x"1fff",x"0000",x"1fff",x"0001",x"0000",x"0001",x"0000",x"1ffd",x"0001",x"0002",x"0000",x"0001",x"0001",x"0000",x"0001",x"0000",x"0000",x"1fff",x"0001",x"0001",x"1ffe",x"1fff",x"1ffe",x"1fff",x"0000",x"0001",x"0001",x"0000",x"1fff",x"1ffe",x"0001",x"0002",x"1fff",x"1ffe",x"0000",x"0000",x"0001",x"0000",x"0000",x"0001",x"0000",x"0003",x"0001",x"0002",x"1ffe",x"0001",x"0001",x"1ffd",x"1fff",x"0001",x"1ffe",x"0000",x"0000",x"1fff",x"0000",x"0000",x"1fff",x"0000",x"0000",x"1ffd",x"1ffe",x"0001",x"0001",x"0002",x"1ffe",x"1fff",x"0000",x"0001",x"1fff",x"0000",x"0001",x"0001",x"0001",x"1fff",x"0000",x"0001",x"0000",x"0002",x"0000",x"0002",x"1ffc",x"0001",x"0000",x"0000",x"0003",x"1ffd",x"0000",x"0002",x"0000",x"1fff",x"0000",x"0000",x"0001",x"1fff",x"0000",x"1fff",x"1fff",x"1fff",x"0001",x"0001",x"1ffd",x"0001",x"1ffe",x"0001",x"1fff",x"0000",x"0002",x"0002",x"1fff",x"1fff",x"1ffe",x"0000",x"0001",x"1ffe",x"0000",x"0001",x"1ffe",x"1fff",x"0000",x"0001",x"0001",x"0003",x"1fff",x"0001",x"0001",x"0002",x"0003",x"1fff",x"0000",x"1fff",x"1fff",x"0001",x"0001",x"1fff",x"0001",x"0000",x"0001",x"0000",x"0000",x"0002",x"0001",x"1ffe",x"0000",x"0001",x"1fff",x"1fff",x"0000",x"1ffe",x"1ffe",x"1ffe",x"0002",x"0001",x"0000",x"0002",x"1fff",x"0000",x"0000",x"0000",x"0000",x"0000",x"0002",x"0001",x"0002",x"1fff",x"1fff",x"1fff",x"1fff",x"1fff",x"1ffe",x"1fff",x"0001",x"1fff",x"1fff",x"0001",
    x"0000",x"0001",x"0001",x"0002",x"0000",x"0002",x"0002",x"0002",x"0002",x"1fff",x"0001",x"0001",x"0002",x"0001",x"0000",x"0002",x"0000",x"1ffe",x"0001",x"1ffe",x"1ffe",x"1ffe",x"0002",x"1fff",x"0001",x"1ffe",x"0000",x"1fff",x"1fff",x"0002",x"0002",x"0001",x"1ffc",x"1fff",x"0002",x"0000",x"0002",x"0000",x"0002",x"0000",x"0002",x"0002",x"1fff",x"0002",x"0000",x"1fff",x"0001",x"0000",x"1ffe",x"1fff",x"1fff",x"0000",x"1fff",x"1fff",x"1fff",x"0000",x"0001",x"1fff",x"0001",x"0001",x"0000",x"0000",x"0002",x"1fff",x"0000",x"0000",x"0002",x"1fff",x"0003",x"1ffe",x"0000",x"1ffd",x"1fff",x"1ffe",x"0001",x"0000",x"0002",x"0002",x"1ffd",x"1ffe",x"1fff",x"0001",x"1fff",x"1ffe",x"1fff",x"1ffe",x"1ffe",x"1ffe",x"0001",x"0001",x"1ffe",x"1ffd",x"1fff",x"0001",x"0002",x"0001",x"0000",x"0002",x"1fff",x"0000",x"0000",x"1fff",x"0002",x"1fff",x"0000",x"0000",x"0001",x"0001",x"0003",x"0002",x"0000",x"0000",x"0002",x"0002",x"1fff",x"1fff",x"1fff",x"0000",x"0001",x"1ffd",x"0001",x"0002",x"0001",x"0000",x"1ffe",x"0001",x"1ffe",x"0000",x"0001",x"0000",x"0000",x"0001",x"0001",x"0002",x"0000",x"0000",x"0000",x"1fff",x"1fff",x"0001",x"0000",x"1fff",x"1ffe",x"0000",x"0000",x"0001",x"1fff",x"1ffe",x"0001",x"0001",x"0002",x"0000",x"0000",x"1ffe",x"1ffe",x"0001",x"0001",x"1fff",x"0001",x"0001",x"0001",x"1fff",x"0001",x"0003",x"0002",x"0002",x"0000",x"1fff",x"0002",x"1ffe",x"0002",x"0001",x"1fff",x"1fff",x"1fff",x"1ffd",x"0001",x"1ffe",x"0000",x"0003",x"0000",x"0003",x"0001",x"1ffe",x"1fff",x"1fff",x"0002",x"1ffe",x"1ffe",x"0001",x"0002",x"0000",x"1ffd",x"0001",x"1ffe",x"0000",x"0001",x"1fff",x"1fff",x"1fff",x"0000",x"1fff",x"1ffe",x"0001",x"0000",x"0002",x"0003",x"0002",x"0000",x"1fff",x"0000",x"1ffe",x"0000",x"1ffd",x"0000",x"1fff",x"1ffd",x"1ffe",x"0001",x"0001",x"1fff",x"1ffe",x"0001",x"1fff",x"0001",x"1ffe",x"0000",x"1fff",x"0001",x"0001",x"1fff",x"0001",x"0002",x"0000",x"0001",x"0000",x"1fff",x"1fff",x"1fff",x"1ffd",x"0001",x"1ffe",x"0001",x"0001",x"0000",x"1fff",x"0000",x"0001",x"1ffe",x"1ffd",x"0001",x"1ffe",x"1fff",x"0002",x"1fff",x"0000",
    x"0001",x"1fff",x"0001",x"0002",x"0001",x"0000",x"0000",x"0000",x"1fff",x"1fff",x"0000",x"0000",x"0000",x"1ffe",x"0000",x"0001",x"0001",x"0001",x"0003",x"0000",x"0001",x"0002",x"1ffd",x"0001",x"1fff",x"0000",x"1fff",x"1ffe",x"0003",x"0003",x"1ffe",x"1ffe",x"1fff",x"1fff",x"1fff",x"0003",x"0001",x"1ffe",x"0001",x"1fff",x"1fff",x"1fff",x"0001",x"1ffe",x"1ffd",x"1fff",x"1ffe",x"1fff",x"1ffd",x"0000",x"0000",x"1ffe",x"0001",x"1ffd",x"1ffe",x"0000",x"0002",x"0000",x"0000",x"1ffe",x"0000",x"1fff",x"0000",x"1ffe",x"1ffe",x"0000",x"1fff",x"0001",x"1ffe",x"0000",x"0001",x"1fff",x"0001",x"0000",x"0000",x"0001",x"1ffe",x"1ffe",x"1ffe",x"0000",x"0002",x"0000",x"0000",x"0000",x"1fff",x"0001",x"0001",x"0001",x"1fff",x"0001",x"0000",x"1ffe",x"1ffd",x"0000",x"1fff",x"0001",x"1fff",x"1fff",x"0001",x"0001",x"0000",x"0002",x"1fff",x"0001",x"0000",x"0002",x"1fff",x"1ffe",x"1ffc",x"0001",x"0000",x"1fff",x"0000",x"1fff",x"1ffe",x"1ffd",x"0001",x"1fff",x"1fff",x"0003",x"1fff",x"1fff",x"1fff",x"0001",x"0001",x"1fff",x"1ffe",x"0001",x"0000",x"0000",x"0001",x"0001",x"0000",x"0000",x"0001",x"1ffe",x"0002",x"0000",x"0000",x"0001",x"0000",x"0000",x"1fff",x"1ffe",x"0000",x"0003",x"0002",x"0000",x"1fff",x"0000",x"0002",x"0000",x"1fff",x"0000",x"0000",x"0000",x"0000",x"0001",x"1fff",x"0002",x"0000",x"0000",x"0001",x"0001",x"0000",x"0001",x"1ffd",x"1ffe",x"1ffe",x"0002",x"0001",x"0001",x"0000",x"0000",x"0000",x"0001",x"1ffd",x"0003",x"0002",x"1fff",x"0000",x"0002",x"0001",x"0002",x"1fff",x"0000",x"0001",x"0000",x"1fff",x"0000",x"1fff",x"1fff",x"1fff",x"1fff",x"1ffe",x"0001",x"1fff",x"0000",x"0000",x"1fff",x"0000",x"0000",x"0001",x"0000",x"1ffe",x"1ffd",x"1fff",x"0001",x"0001",x"0000",x"0001",x"1ffe",x"1fff",x"0002",x"0000",x"1fff",x"0000",x"0002",x"0000",x"0000",x"1fff",x"1ffe",x"1fff",x"0000",x"1fff",x"0000",x"1fff",x"0001",x"0000",x"0000",x"0002",x"1ffe",x"0001",x"0000",x"0003",x"0000",x"0002",x"0002",x"0000",x"0000",x"0000",x"0001",x"0002",x"0000",x"0000",x"1ffe",x"0000",x"1ffe",x"1fff",x"0002",x"1fff",x"0000",x"0000",x"0003",x"0001",x"1ffd",    
    --pkh
    x"4937", x"6c18", x"232e", x"98d7", x"b2e7", x"80aa", x"e42a", x"2615", x"21d7", x"ed7d", x"0ac7", x"59fc", x"ca99", x"9d89", x"580a", x"f660", 
    
      --z
    x"aca6", x"7585", x"16a0", x"42ca", x"e90d", x"9212", x"2afa", x"109c", x"9357", x"8213", x"c92f", x"62e0", x"a9a5", x"d85e", x"10bc", x"4bc1", 
    
    --SK--share1=======================================================================================================
--    --S polyvec 
--    x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
--    x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
--    x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
--    x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
--    x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
--    x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
--    x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
--    x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
    
--    x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
--    x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
--    x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
--    x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
--    x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
--    x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
--    x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
--    x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
    
--    x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
--    x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
--    x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
--    x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
--    x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
--    x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
--    x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
--    x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
    -- randmoly shared S polyvec
    
    x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
    x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
    x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
    --rand shared
 
    --PKH
    x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
    x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
   
    --Z
    x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
    x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",

    --cipher = (Bp, cm)=========================================================
    --Bp
   --cipher = (Bp, cm)=========================================================
    --Bp

    x"4b91", x"0f96", x"a773", x"9880", x"9dc6", x"2bc4", x"7e75", x"143b", x"7711", x"c245", x"2ef3", x"e627", x"42e6", x"cb0c", x"14f0", x"3afb", x"a334", x"61b5", x"46d9", x"7461", x"d5d1", x"4b24", x"0f15", x"6ac4", x"52a5", x"09cb", x"1d9a", x"0b0d", x"5641", x"241c", x"38af", x"186e", x"b94e", x"0e13", x"b08d", x"5e0f", x"f855", x"7288", x"6f0e", x"c455", x"5228", x"7bed", x"c205", x"de7e", x"bfc6", x"70a6", x"fc2d", x"d37f", x"9ba9", x"7730", x"557b", x"6203", x"32c6", x"b999", x"d60c", x"7df1", x"941c", x"0a9e", x"3cc2", x"94de", x"ae67", x"8f6b", x"f06c", x"19ea", x"9b1f", x"5ce7", x"31ea", x"9806", x"e5c3", x"dab1", x"ec28", x"427e", x"f01f", x"66fd", x"64fe", x"52eb", x"0cfc", x"d721", x"3738", x"f791", x"5091", x"e8d1", x"42b3", x"2b35", x"be60", x"36f2", x"c7e8", x"a619", x"3f68", x"035a", x"7c57", x"15ff", x"fa6d", x"28e3", x"23ed", x"72ed", x"a2bb", x"400c", x"a3c3", x"bd67", x"3051", x"68e7", x"0ad6", x"9c0c", x"e8fb", x"c393", x"cfa4", x"efa2", x"d5a1", x"0116", x"9e0c", x"628f", x"66c4", x"25ef", x"6418", x"830a", x"d3e8", x"7813", x"5f95", x"95a7", x"f9e8", x"7156", x"0f03", x"0cef", x"b8b0", x"b3b7", x"438f", x"919a", x"4247", x"4ca8", x"ee15", x"170c", x"b158", x"30bd", x"e3c5", x"d380", x"a645", x"fc7d", x"11d5", x"4d6b", x"63a2", x"e654", x"5885", x"7851", x"9650", x"8e40", x"9be9", x"1e61", x"fd5c", x"6902", x"3286", x"1b41", x"80ac", x"a7fc", x"271e", x"0f51", x"763c", x"8a51", x"b467", x"b23e", 

    x"5b51", x"e5e4", x"1d16", x"4680", x"ba16", x"1a51", x"c613", x"ca95", x"e098", x"0454", x"7b28", x"2a8f", x"4a99", x"9dda", x"1e89", x"1959", x"1ecd", x"ffad", x"9e8a", x"a8bd", x"6d3b", x"e845", x"12d0", x"c0d0", x"e45d", x"aa95", x"1181", x"c898", x"81bd", x"4c8b", x"cf64", x"2006", x"363f", x"a7f6", x"e297", x"84da", x"f7d5", x"56b3", x"7ded", x"d604", x"e9bf", x"408f", x"7a14", x"6996", x"e2a8", x"271e", x"7b38", x"fa9e", x"cd75", x"d83e", x"97a6", x"4918", x"f4a9", x"6802", x"52ee", x"73c6", x"0172", x"eeb8", x"97b2", x"24a5", x"82b6", x"2d84", x"1a05", x"d8d1", x"8848", x"4dd0", x"d3fd", x"5fd5", x"8e98", x"c147", x"acb0", x"84ed", x"08b2", x"6385", x"1f5d", x"0c2f", x"fd59", x"8506", x"ea6b", x"f327", x"dc4b", x"d2a1", x"1915", x"1288", x"62e6", x"f880", x"af42", x"7792", x"4d1b", x"94f2", x"6054", x"1e82", x"084b", x"1fc1", x"b783", x"a60f", x"777c", x"1bdc", x"4fe1", x"33ef", x"f08f", x"6edf", x"e6dd", x"2f68", x"0af0", x"a19d", x"6115", x"40f7", x"2345", x"f444", x"3c36", x"7ca0", x"49c8", x"13a5", x"2d93", x"41e9", x"2005", x"74c6", x"288f", x"5835", x"19cc", x"b38a", x"0a89", x"28c2", x"1e0a", x"fa62", x"0b5c", x"fab2", x"8270", x"4391", x"7004", x"f51e", x"ad92", x"a1a1", x"9c31", x"8a47", x"8987", x"a101", x"b6da", x"c09a", x"4820", x"530e", x"771a", x"de1b", x"9332", x"c8c7", x"491f", x"d6e9", x"c2b7", x"0247", x"3f2b", x"ec1f", x"6f0d", x"38d8", x"8592", x"f564", x"8ce8", x"76f8", x"2bbd", x"c04e", 

    x"485c", x"cef1", x"47fb", x"6bcb", x"ac1e", x"7863", x"67d0", x"ea41", x"b2f9", x"bc09", x"b0c5", x"3b5f", x"29de", x"6bdf", x"368d", x"8b41", x"be11", x"0922", x"5573", x"d198", x"d3f2", x"24e0", x"6ef5", x"6581", x"7053", x"716f", x"b251", x"7a7b", x"a53a", x"da7d", x"07e7", x"7060", x"3d0d", x"2793", x"57b8", x"ec8b", x"1767", x"e7c7", x"59e8", x"87d1", x"75a8", x"1d98", x"19d3", x"1edc", x"d4e4", x"de7f", x"d294", x"26ca", x"f01a", x"ede3", x"590d", x"4938", x"371d", x"d615", x"abee", x"f5f8", x"10e9", x"7870", x"ff94", x"5f25", x"1bff", x"9113", x"6667", x"01a0", x"5e39", x"5dc1", x"fbc1", x"10c9", x"dc2a", x"c169", x"04c3", x"3c47", x"d412", x"0d67", x"5a0c", x"3b8e", x"41e5", x"4b90", x"8c95", x"7ff0", x"2adc", x"4e92", x"9364", x"c769", x"4274", x"2970", x"7edd", x"8057", x"10a7", x"3e2e", x"0093", x"08e0", x"7e75", x"46f1", x"e203", x"6288", x"b9c3", x"0eb0", x"d401", x"e49c", x"6501", x"81a3", x"8c5f", x"f013", x"30bf", x"77da", x"64a4", x"c7c8", x"e19c", x"ea5b", x"faf7", x"5f95", x"f722", x"4bbb", x"9873", x"16b9", x"d57f", x"8171", x"d167", x"9732", x"f3db", x"8085", x"e8a2", x"ae2e", x"1631", x"141c", x"fe53", x"ed08", x"d12f", x"d0fa", x"9678", x"db34", x"4aea", x"3c56", x"e53a", x"fdaa", x"6547", x"d3ef", x"1e44", x"ac47", x"1429", x"deef", x"019e", x"c2cf", x"a919", x"b079", x"7511", x"2a29", x"8509", x"2742", x"b627", x"d38a", x"cd13", x"315b", x"a437", x"40ec", x"e6fb", x"d3bb", x"85f2", x"f907", 
    
    --cm
    x"44d0", x"a9c5", x"1054", x"2e34", x"2132", x"bf4c", x"6713", x"1fc3", x"55ce", x"bf6c", x"1853", x"8f99", x"9b67", x"5619", x"628e", x"c315", x"59b3", x"8ab3", x"7fc7", x"9cfa", x"31ff", x"3f61", x"4740", x"9d88", x"c103", x"34b7", x"cfb4", x"aefb", x"75b3", x"c3bd", x"4059", x"bbd8", x"8eff", x"1e03", x"2eeb", x"16c6", x"738c", x"4079", x"9e97", x"2deb", x"be28", x"e948", x"8545", x"5866", x"30b2", x"56f9", x"977e", x"6853", x"9620", x"8f84", x"e5f7", x"3c35", x"119c", x"63db", x"a33e", x"c38d", x"eb79", x"0448", x"9abf", x"3242", x"e5ce", x"5636", x"2acb", x"c4d2", 
    --end chipertext
    --end chipertext
    
    others=>x"0000"
    );
    

end decaps_tv_shared_pkg_2;

package body decaps_tv_shared_pkg_2 is
end package body;
