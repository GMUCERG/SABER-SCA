--------------------------------------------------------------------------------
--! @file       decaps_tv_shared_pkg.vhd
--! @author     Abubakr Abdulgadir
--! @copyright  Copyright (c) 2021 Cryptographic Engineering Research Group
--!             ECE Department, George Mason University Fairfax, VA, U.S.A.
--!             All rights Reserved.
--------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.all;
use ieee.numeric_std.all;

use work.saber_pkg.all;
use work.saber_pr_pkg.all;

package decaps_tv_shared_pkg is


    type decaps_input_shared_arr_type is array (0 to 2**DIN_FIFO_LOG2DEPTH-1) of std_logic_vector(DIN_FIFO_WIDTH-1 downto 0);
    constant DECAPS_INPUT_DATA : decaps_input_shared_arr_type := 
    (
    --opcode =================================================================================================
    OPCODE_DECAPS,
    --PK======================================================================================================
    --b polycev
    x"aeeb", x"17a9", x"b67a", x"db0c", x"e521", x"dfb6", x"9f96", x"af19", x"0773", x"a31f", x"0b05", x"a84c", 
    x"7e90", x"fe9b", x"5a38", x"e4e7", x"f1e9", x"4ab6", x"3bbf", x"8306", x"9d61", x"4612", x"a7d3", x"ce24", 
    x"932c", x"b5c4", x"6277", x"59d8", x"be47", x"89a2", x"4269", x"aae8", x"7b1e", x"f3b2", x"baff", x"a251", 
    x"d996", x"917f", x"c333", x"c7a8", x"fd4d", x"e318", x"e58d", x"24b5", x"410e", x"85e8", x"6891", x"8405", 
    x"c624", x"df5c", x"d19c", x"5290", x"f802", x"5a8a", x"72f7", x"851f", x"4106", x"f274", x"27f9", x"7db9", 
    x"8169", x"5fce", x"1f26", x"1fa2", x"befa", x"bb74", x"793b", x"23b3", x"48a5", x"a722", x"a605", x"81a6", 
    x"c257", x"d1ee", x"7af3", x"5c9f", x"a169", x"a6d5", x"c167", x"35ba", x"bfd4", x"f16f", x"1fd2", x"bb37", 
    x"0e09", x"5593", x"eedd", x"3a4b", x"a887", x"e8cc", x"a138", x"a7b0", x"a7f6", x"5147", x"484b", x"08b2", 
    x"d398", x"af64", x"a1cc", x"dc32", x"520f", x"12fb", x"3c07", x"5d23", x"1f28", x"037b", x"1b34", x"1b0a", 
    x"a60b", x"64ee", x"d6dc", x"41d6", x"3d38", x"4782", x"881e", x"6a2a", x"9f95", x"a88e", x"7542", x"a557", 
    x"f0a3", x"65ee", x"f005", x"d5d4", x"992c", x"1f05", x"feb6", x"a9c2", x"734e", x"8361", x"2667", x"a9b8", 
    x"f427", x"a858", x"189d", x"58d0", x"9e9f", x"fbc2", x"1928", x"57e1", x"976f", x"ec72", x"620b", x"298c", 
    x"7de8", x"35fc", x"a2ed", x"ba6a", x"d51d", x"a966", x"6dca", x"05ba", x"9c51", x"cfcd", x"0964", x"5b22", 
    x"7618", x"3f15", x"ca43", x"2d0b", x"96ef", x"a597", x"3aa5", x"9b44", x"e146", x"a7ea", x"3fbc", x"4e05", 
    x"a85d", x"b63a", x"088c", x"a06e", x"a9c9", x"328c", x"6529", x"b4e9", x"6d46", x"c652", x"831b", x"23c6", 
    x"ee45", x"8ba2", x"4ce1", x"c9b5", x"456f", x"1e47", x"eff7", x"7660", x"e3af", x"3fdf", x"a8a7", x"9988", 
    x"2ec6", x"bf32", x"bfdc", x"88df", x"6497", x"1345", x"8c80", x"a210", x"bf09", x"38fa", x"eaf7", x"e694", 
    x"0fac", x"9b13", x"b8c3", x"ffad", x"afc4", x"7436", x"3056", x"3dbe", x"50a7", x"7738", x"977e", x"fe9c", 
    x"c4c0", x"19bd", x"0e47", x"dc1c", x"292f", x"dc86", x"42b2", x"70fb", x"567f", x"2e33", x"3b75", x"b90d", 
    x"688e", x"08c1", x"8797", x"f1c2", x"b3db", x"8e3f", x"1c02", x"8952", x"44d6", x"650d", x"2761", x"e64f", 
    x"14ff", x"0186", x"c9bf", x"3a39", x"501a", x"dfa9", x"111a", x"74a2", x"8047", x"f06b", x"1249", x"c2e9", 
    x"3c10", x"e735", x"8eba", x"43c9", x"b432", x"aeda", x"d7a0", x"9a9f", x"ad21", x"457e", x"5709", x"46b1", 
    x"3b8d", x"47a4", x"e677", x"4f5e", x"b434", x"8010", x"90ce", x"3b0d", x"46cb", x"69eb", x"a271", x"4651", 
    x"5bbd", x"1da9", x"ac0c", x"c8e1", x"3b30", x"1062", x"bcf1", x"49e6", x"fdcc", x"ed92", x"6110", x"8ace", 
    x"8f46", x"89e6", x"e5c8", x"e2de", x"2d8c", x"f75c", x"881a", x"b3c1", x"42fd", x"0382", x"979b", x"0d29", 
    x"23e9", x"5adc", x"e002", x"1cce", x"6e6f", x"54af", x"4b50", x"7a22", x"1844", x"193c", x"794a", x"f59c", 
    x"fb70", x"7d01", x"526a", x"88bb", x"f8df", x"c062", x"b3fd", x"df17", x"5bdb", x"4c3a", x"9a57", x"0099", 
    x"4723", x"a005", x"87cd", x"6a8a", x"f123", x"06e9", x"cb4b", x"8e15", x"d792", x"68e4", x"5f75", x"e93c", 
    x"2c6d", x"24d9", x"930e", x"6be9", x"c6ef", x"4273", x"6f23", x"b74b", x"54fe", x"a535", x"f092", x"6d95", 
    x"70f2", x"89d9", x"1cc2", x"6309", x"c65e", x"c95a", x"fbb2", x"ad42", x"d6ab", x"89a4", x"a8e3", x"fbad", 
    x"3bf1", x"5ec5", x"7e96", x"ba72", x"cda5", x"85cc", x"f504", x"5ead", x"80e1", x"ffcc", x"8f56", x"bc0c", 
    x"33cf", x"fe02", x"90d2", x"45db", x"ad11", x"1281", x"cf69", x"ec41", x"ae9c", x"5b0e", x"b192", x"f154", 
    x"d5c6", x"38d2", x"f64d", x"cf29", x"00aa", x"c0da", x"7e54", x"d32f", x"fe7c", x"dae3", x"d5d7", x"33a0", 
    x"37f6", x"cdcc", x"53ae", x"e04d", x"e609", x"2a92", x"873d", x"17d6", x"6676", x"5246", x"5c88", x"5ea5", 
    x"9ab3", x"bbab", x"ecab", x"a966", x"71cd", x"2d82", x"5f48", x"c03d", x"f6a0", x"68dd", x"2559", x"26bf", 
    x"e434", x"5388", x"2cc2", x"7cc0", x"1ab1", x"5e3f", x"3db9", x"db07", x"84b9", x"6397", x"0134", x"eae8", 
    x"0716", x"3fb0", x"770c", x"03d8", x"7eef", x"fd61", x"1f22", x"b2c0", x"853a", x"2436", x"2fd9", x"d695", 
    x"5e06", x"b278", x"47ec", x"90ac", x"c123", x"c0dc", x"276b", x"9ec9", x"4960", x"feb5", x"f667", x"914b", 
    x"e730", x"7641", x"185c", x"a9ad", x"f7be", x"6f29", x"eb4a", x"745c", x"195e", x"a94c", x"bb2d", x"02d6", 
    x"f4f0", x"c636", x"f10c", x"e6e8", x"012d", x"5ef9", x"9fcd", x"a0cb", x"6f4f", x"b53c", x"bfc1", x"397e", 
    --SEED_A
    x"8807", x"a700", x"66a7", x"5ebe", x"4a24", x"fcd3", x"9ee2", x"8339", x"fe9c", x"c982", x"abaa", x"7cf2", 
    x"2fcf", x"53c6", x"2d56", x"8f93",
    --SEED_A second share (no need to share but this is just a work around since SHA3 needs 2 shares).
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000",
    --END_PK===================================================================================================
    
    --SK--share0=======================================================================================================
    --S polyvec 
       --orig
--    x"0001",x"1fff",x"0000",x"0000",x"1ffe",x"0002",x"0001",x"0000",x"1fff",x"0001",x"0000",x"0001",x"1ffe",x"1fff",x"0003",x"1fff",x"1ffe",x"1ffd",x"1fff",x"0003",x"0001",x"0002",x"0000",x"0001",x"0002",x"0002",x"1fff",x"0000",x"0000",x"1fff",x"0001",x"0000",x"1ffe",x"0000",x"1ffc",x"0000",x"0001",x"0000",x"1fff",x"0000",x"1fff",x"0001",x"0000",x"1ffe",x"1ffd",x"0000",x"1ffe",x"1ffd",x"1fff",x"1fff",x"1fff",x"0000",x"1fff",x"1fff",x"1ffe",x"0001",x"0000",x"0000",x"1fff",x"1fff",x"0000",x"0001",x"0001",x"0002",x"0000",x"0001",x"0001",x"0002",x"1fff",x"0000",x"0000",x"0000",x"0001",x"0001",x"0001",x"0003",x"0001",x"0001",x"1fff",x"1fff",x"1ffd",x"0001",x"1fff",x"0001",x"1fff",x"0000",x"1ffe",x"0001",x"1fff",x"0001",x"1ffe",x"0000",x"1ffe",x"1ffe",x"0001",x"0000",x"0000",x"0000",x"0000",x"0001",x"0001",x"1fff",x"1fff",x"0000",x"0001",x"0000",x"1fff",x"0001",x"0001",x"1ffd",x"1ffe",x"0000",x"0003",x"1ffe",x"0000",x"0002",x"1ffe",x"0000",x"0001",x"0003",x"0000",x"0001",x"0001",x"0001",x"1fff",x"1ffd",x"1ffe",x"0000",x"1ffe",x"0000",x"0001",x"1fff",x"1fff",x"1ffe",x"0001",x"0000",x"1fff",x"0002",x"1fff",x"0000",x"0004",x"0001",x"1ffe",x"0003",x"1fff",x"0002",x"0001",x"0002",x"0003",x"0000",x"1fff",x"0000",x"0000",x"1ffe",x"1fff",x"0000",x"1fff",x"0000",x"0002",x"1fff",x"0001",x"0001",x"1ffe",x"1fff",x"1ffd",x"0000",x"0002",x"0000",x"0002",x"0000",x"0002",x"0001",x"1ffe",x"1fff",x"1ffe",x"0000",x"0000",x"1fff",x"0003",x"1ffe",x"0000",x"0000",x"1ffe",x"0001",x"0001",x"0001",x"0001",x"0000",x"0000",x"0000",x"0002",x"1fff",x"1fff",x"0001",x"0000",x"0001",x"1fff",x"0001",x"0000",x"0001",x"1ffd",x"1ffe",x"0000",x"0000",x"1ffe",x"1fff",x"1fff",x"0000",x"0001",x"0001",x"1fff",x"0001",x"0001",x"0002",x"1ffe",x"1ffe",x"0001",x"1ffe",x"0002",x"0000",x"1ffe",x"0001",x"1fff",x"0000",x"1fff",x"1fff",x"0001",x"1fff",x"1ffe",x"0002",x"1ffe",x"0001",x"0001",x"0000",x"0000",x"1fff",x"0000",x"1fff",x"1fff",x"0001",x"0002",x"0001",x"1fff",x"0000",x"0001",x"0002",x"1fff",x"0001",x"0002",x"0001",x"0001",x"1fff",x"0000",x"0000",x"1fff",x"0001",
--    x"1fff",x"0000",x"0000",x"0001",x"1fff",x"0000",x"0000",x"0001",x"0003",x"1fff",x"0001",x"0000",x"0001",x"0000",x"1ffe",x"0001",x"0001",x"0001",x"1ffe",x"1fff",x"0002",x"1fff",x"1ffd",x"0001",x"1fff",x"0001",x"0000",x"0000",x"0001",x"0003",x"1ffe",x"1ffd",x"0000",x"0000",x"0000",x"1fff",x"0000",x"1ffe",x"0000",x"0001",x"0000",x"0000",x"0000",x"0000",x"0001",x"0002",x"0000",x"0001",x"1ffd",x"0000",x"1fff",x"0002",x"1ffe",x"1ffe",x"0002",x"0001",x"0001",x"0002",x"0002",x"0000",x"1ffe",x"0000",x"0000",x"1ffe",x"0001",x"0001",x"0001",x"0002",x"0001",x"0001",x"0001",x"1ffe",x"0000",x"0001",x"0002",x"1fff",x"0002",x"0002",x"1fff",x"1fff",x"1fff",x"0003",x"0000",x"0000",x"1ffe",x"0001",x"0000",x"0000",x"0000",x"0001",x"0000",x"0001",x"0000",x"1fff",x"1fff",x"0000",x"0001",x"0001",x"1fff",x"1fff",x"0000",x"1ffe",x"0002",x"1fff",x"1ffe",x"0000",x"1fff",x"0002",x"0002",x"0000",x"0000",x"0000",x"0000",x"0000",x"1fff",x"0000",x"0000",x"0001",x"0000",x"1fff",x"0000",x"0000",x"0002",x"0001",x"0001",x"1fff",x"0001",x"0001",x"0000",x"0003",x"1fff",x"0001",x"0003",x"1fff",x"1fff",x"0002",x"0000",x"0000",x"0001",x"0000",x"1fff",x"0003",x"0000",x"1ffe",x"1ffe",x"0000",x"1ffe",x"0002",x"0001",x"1ffd",x"0002",x"0001",x"0001",x"1fff",x"0000",x"0000",x"0000",x"1fff",x"0001",x"0001",x"1ffe",x"0002",x"0002",x"1fff",x"0003",x"0001",x"0000",x"0000",x"0002",x"0001",x"0001",x"1ffe",x"1fff",x"0001",x"0001",x"0000",x"0000",x"1fff",x"0001",x"1fff",x"1ffd",x"0002",x"1fff",x"1ffe",x"1fff",x"1ffe",x"0001",x"1ffd",x"0001",x"0001",x"0002",x"0000",x"0001",x"0001",x"0000",x"0000",x"0001",x"1fff",x"1fff",x"1fff",x"0001",x"0001",x"0000",x"0003",x"0001",x"0000",x"0000",x"0000",x"1fff",x"0000",x"0002",x"1fff",x"1ffe",x"0001",x"1fff",x"0002",x"0000",x"0002",x"0002",x"0001",x"0001",x"1ffd",x"0000",x"0001",x"0000",x"0000",x"0000",x"0002",x"0000",x"0001",x"0001",x"0002",x"0000",x"0000",x"0001",x"0001",x"0000",x"1fff",x"1fff",x"0001",x"0000",x"0002",x"1ffe",x"0004",x"1fff",x"1ffe",x"1fff",x"1ffe",x"0000",x"1fff",x"0002",x"0001",x"0001",x"1fff",x"0000",x"1ffe",
--    x"1ffe",x"0000",x"0002",x"1fff",x"0000",x"1ffe",x"1ffe",x"1ffe",x"0000",x"0002",x"0000",x"1fff",x"1fff",x"1fff",x"0001",x"0000",x"0002",x"0003",x"0000",x"1ffe",x"0001",x"1ffd",x"0002",x"0002",x"0001",x"0001",x"1fff",x"1fff",x"1fff",x"0000",x"0000",x"0000",x"0000",x"0000",x"0001",x"0001",x"0001",x"1ffe",x"1ffe",x"1fff",x"0000",x"0002",x"1ffd",x"0001",x"0000",x"0001",x"0001",x"0001",x"1fff",x"1fff",x"0001",x"1ffd",x"0002",x"1fff",x"1fff",x"1ffe",x"1fff",x"0002",x"0000",x"1ffe",x"0001",x"0001",x"1fff",x"0001",x"1ffc",x"1fff",x"0001",x"0002",x"0001",x"0000",x"0000",x"1fff",x"0001",x"0000",x"0001",x"0000",x"1ffe",x"0001",x"1ffd",x"0001",x"0001",x"0000",x"1fff",x"1ffe",x"0001",x"1fff",x"0002",x"1fff",x"1ffe",x"0000",x"0002",x"1ffe",x"0000",x"1fff",x"0000",x"0001",x"0001",x"1ffc",x"0002",x"1fff",x"1ffe",x"0001",x"0001",x"0001",x"0001",x"0000",x"1fff",x"1fff",x"0000",x"1fff",x"1ffe",x"0000",x"1ffe",x"0001",x"0003",x"0000",x"1ffe",x"0002",x"0000",x"1fff",x"0000",x"1fff",x"0000",x"1fff",x"1ffe",x"0002",x"1ffe",x"1fff",x"1fff",x"0002",x"1ffe",x"0000",x"1ffd",x"1fff",x"0000",x"1ffd",x"0001",x"0001",x"1fff",x"1fff",x"0000",x"0000",x"1fff",x"1ffe",x"1ffe",x"0001",x"1ffd",x"0001",x"1ffe",x"1ffe",x"1fff",x"1fff",x"0001",x"1fff",x"0000",x"0001",x"0000",x"0000",x"0000",x"1fff",x"0000",x"0001",x"0002",x"0001",x"1fff",x"0003",x"0001",x"0001",x"0001",x"0001",x"1ffe",x"0000",x"1ffe",x"1fff",x"0000",x"1ffe",x"1ffe",x"1fff",x"1fff",x"1fff",x"0001",x"0000",x"0001",x"1fff",x"0001",x"0001",x"0001",x"0000",x"1fff",x"0000",x"0001",x"0001",x"1fff",x"0001",x"1fff",x"0002",x"0001",x"0002",x"0000",x"0001",x"1ffe",x"0001",x"0001",x"0000",x"0001",x"0001",x"0000",x"1ffe",x"0002",x"0001",x"0000",x"0002",x"0003",x"1fff",x"0001",x"0000",x"0000",x"0001",x"0001",x"0001",x"0001",x"0000",x"0002",x"0000",x"1fff",x"0001",x"1ffe",x"0002",x"0001",x"1fff",x"0000",x"0001",x"0000",x"1ffe",x"1fff",x"1fff",x"1ffe",x"1ffe",x"1fff",x"1ffe",x"0002",x"0000",x"1fff",x"1ffe",x"0000",x"1ffe",x"1fff",x"0001",x"1fff",x"1fff",x"0001",x"0000",x"1fff",x"1ffe",x"0001",x"0002",
    --rand shared
    x"1f53",x"1ede",x"17cd",x"1587",x"0cd3",x"18e3",x"1135",x"01f5",x"0d3e",x"159d",x"02d4",x"0e08",x"13ca",x"0329",x"13a2",x"04ae",x"1bbd",x"0acb",x"0cfd",x"02c8",x"1675",x"0537",x"1fd5",x"06f4",x"1a44",x"012f",x"0a07",x"00f8",x"1138",x"1055",x"0456",x"1d46",x"0013",x"0eab",x"1546",x"1560",x"0dfb",x"1165",x"0556",x"0969",x"1f15",x"06f4",x"1c8b",x"14ab",x"1043",x"16e0",x"139d",x"0b95",x"04d1",x"1d45",x"0eef",x"09db",x"1901",x"0aa1",x"0da8",x"156b",x"1467",x"0af9",x"06ab",x"0833",x"0be5",x"1d5e",x"01d2",x"09b6",x"07cf",x"0efc",x"1133",x"09ad",x"04e8",x"0d5d",x"0084",x"0ab8",x"1db0",x"1778",x"01ea",x"1994",x"0310",x"0435",x"07d5",x"02c2",x"1594",x"0fed",x"03b8",x"1198",x"1f2b",x"1d54",x"02ed",x"16bf",x"040f",x"0d61",x"1918",x"0d58",x"0968",x"1e5b",x"1d3d",x"1283",x"0993",x"028c",x"1072",x"0d2c",x"074a",x"1989",x"0abf",x"03dc",x"1175",x"1eae",x"06df",x"1dd7",x"1f8d",x"1e45",x"1ead",x"07e8",x"1c87",x"0529",x"026e",x"0190",x"14b2",x"1b27",x"0823",x"076a",x"191c",x"0675",x"0451",x"0825",x"1201",x"19d1",x"191e",x"1c22",x"1f74",x"1403",x"1da1",x"08ab",x"0d59",x"0601",x"0162",x"1db8",x"1731",x"1c67",x"1328",x"0c52",x"0229",x"0136",x"1bd5",x"06af",x"065c",x"077f",x"1fc1",x"0b29",x"0f26",x"158c",x"08cf",x"139c",x"1519",x"18fb",x"04f2",x"0035",x"1dd6",x"1ebf",x"1d5b",x"044d",x"06a1",x"09ce",x"0975",x"0388",x"1cc4",x"082e",x"0e76",x"1355",x"1ead",x"1ddc",x"1716",x"010e",x"0900",x"11b2",x"01e5",x"08b6",x"14b2",x"0b89",x"0721",x"0cf4",x"0628",x"02a8",x"1af3",x"0787",x"039a",x"0e9d",x"07b2",x"10b9",x"0611",x"027e",x"190a",x"092b",x"1bbe",x"10e1",x"1fc1",x"12e6",x"0f7d",x"1313",x"0cdd",x"1186",x"1c05",x"0cc4",x"05c2",x"1ef7",x"0da8",x"09e8",x"0fd0",x"1347",x"17a8",x"0b18",x"04d7",x"16b4",x"0d7a",x"1a96",x"1629",x"1306",x"1878",x"1cce",x"0233",x"02a7",x"1bff",x"1218",x"1c1f",x"0e94",x"1e92",x"1323",x"1de0",x"1ad4",x"1458",x"19e0",x"165b",x"1f2c",x"1ffa",x"0364",x"15d2",x"1096",x"05e2",x"139f",x"1eb2",x"1f12",x"09fc",x"0c4e",x"0e07",x"020b",x"06bf",x"16ca",x"1bb9",x"153a",x"0a26",x"04a9",x"1bd6",x"1fc0",x"0422",x"00d1",x"11aa",x"1fb4",x"0c46",x"0c83",x"1ba8",x"1f7b",x"105b",x"0bcc",x"06a7",x"00d5",x"1319",x"1f00",x"106b",x"0fa2",x"057d",x"1bc1",x"1770",x"0a2b",x"0aa5",x"0fee",x"106b",x"05d9",x"13d7",x"0f2a",x"0df3",x"02c4",x"0eb4",x"01c7",x"145d",x"1801",x"1017",x"18d7",x"0158",x"1959",x"1945",x"1796",x"1ff1",x"1450",x"195f",x"0cf0",x"06c0",x"11f2",x"07c3",x"0161",x"0f1f",x"15c6",x"1434",x"1e40",x"1708",x"1b18",x"1446",x"054b",x"0fc4",x"0f3e",x"04f5",x"0465",x"0f47",x"05f7",x"0619",x"09b3",x"0b2a",x"1a85",x"0fa5",x"1384",x"02fc",x"16ff",x"0bbe",x"072a",x"1bf9",x"0c0c",x"0b10",x"1cb9",x"1e45",x"000d",x"070b",x"0fd6",x"096a",x"1d27",x"1500",x"0198",x"0b70",x"1a9b",x"0377",x"0a9e",x"14d8",x"1bdc",x"0598",x"16ff",x"0b7e",x"145e",x"0a79",x"17b4",x"016e",x"1aa0",x"1fbe",x"1f3d",x"15ee",x"03e3",x"0c56",x"1b2f",x"1288",x"1e03",x"0264",x"1ab4",x"18ce",x"173c",x"16e4",x"033b",x"05d1",x"03bb",x"17d3",x"0558",x"0858",x"1063",x"14f2",x"0f41",x"00cc",x"1954",x"1c07",x"0456",x"172c",x"12f8",x"10cf",x"0c20",x"1421",x"0d4d",x"0681",x"0e03",x"01a7",x"00f8",x"05be",x"003e",x"0e64",x"1be6",x"091b",x"13ba",x"1662",x"056d",x"10e6",x"0daf",x"0799",x"0550",x"0cf0",x"0c72",x"15ff",x"1cc9",x"0a99",x"0dc0",x"170f",x"1df5",x"0450",x"1eea",x"19fd",x"1664",x"0007",x"0d97",x"04f1",x"1928",x"0226",x"1f6d",x"0a25",x"0671",x"0665",x"05c4",x"0ce2",x"0f56",x"0fbc",x"0cfa",x"0d31",x"121e",x"0efb",x"16e1",x"15db",x"0d47",x"1ecd",x"06d9",x"05a5",x"079f",x"12e4",x"04fa",x"0bb1",x"07af",x"1935",x"0267",x"0688",x"0712",x"1bd4",x"1c19",x"01a7",x"07dd",x"1102",x"0de8",x"16b2",x"14d1",x"0268",x"0e67",x"1261",x"1403",x"181a",x"11b5",x"0c6f",x"07d8",x"08bf",x"04ff",x"1fff",x"1171",x"11de",x"1273",x"01b9",x"1441",x"1e6a",x"0352",x"1947",x"16ab",x"0a45",x"1b3a",x"19a8",x"0665",x"1693",x"0c22",x"0cd5",x"0be4",x"1858",x"025e",x"0ec1",x"1280",x"10d8",x"016d",x"172f",x"1b78",x"0204",x"0840",x"05a4",x"0e3c",x"0eb2",x"0cb7",x"01d4",x"1f44",x"1705",x"16bd",x"0dce",x"0416",x"1fcf",x"1053",x"134c",x"193d",x"18a7",x"0b20",x"1eb9",x"0c1e",x"1d54",x"0194",x"09ba",x"0245",x"11ca",x"1158",x"1ccb",x"1b95",x"08fc",x"1946",x"02c1",x"0db4",x"120d",x"1f4f",x"1e6f",x"1f2b",x"17d5",x"0343",x"18dd",x"0409",x"0236",x"1358",x"0ab7",x"19e4",x"0bfc",x"167a",x"0337",x"10b8",x"0d31",x"1914",x"1da5",x"0fb5",x"1f3d",x"0fee",x"05d3",x"0f28",x"057e",x"1243",x"1125",x"1683",x"1dd4",x"0ba6",x"12de",x"1b21",x"1459",x"1ca9",x"1eec",x"0df7",x"1016",x"15e5",x"0942",x"0239",x"0e9b",x"11ee",x"00f3",x"1ce5",x"0c3a",x"0478",x"089c",x"03bc",x"08e3",x"0b2f",x"1521",x"1b99",x"1e76",x"19ca",x"10e7",x"15c8",x"05d1",x"0cd9",x"0307",x"0fb3",x"051d",x"18a7",x"01a9",x"1f14",x"0521",x"1671",x"0078",x"04fc",x"160a",x"1e4c",x"162f",x"0582",x"02e0",x"13d8",x"1135",x"1545",x"0993",x"1580",x"0991",x"01d7",x"0e6e",x"1bd4",x"003a",x"0be4",x"1ea4",x"058c",x"06ac",x"16e4",x"0b4f",x"19a5",x"0076",x"1198",x"06ad",x"00b4",x"0f54",x"037a",x"1abc",x"0187",x"076e",x"0417",x"1b14",x"0845",x"1907",x"0324",x"1c6f",x"1689",x"14c5",x"1519",x"1221",x"15d4",x"0a40",x"08a1",x"0c53",x"1dc9",x"1102",x"1610",x"0c7e",x"0c57",x"073d",x"0f3a",x"1672",x"0c19",x"107a",x"0baa",x"02d0",x"1391",x"0028",x"1d3c",x"1d51",x"0dfa",x"1cfd",x"11f1",x"16e5",x"01a9",x"05a6",x"0ccc",x"04c6",x"016f",x"0518",x"0d21",x"19ce",x"10c5",x"1409",x"0025",x"1566",x"178b",x"0399",x"0710",x"1c53",x"1f3d",x"0d7a",x"0797",x"05b2",x"1279",x"1770",x"0e09",x"172a",x"19a9",x"06e9",x"0be7",x"181a",x"1d77",x"0276",x"032a",x"183e",x"070b",x"1bc7",x"0bdb",x"04a0",x"127d",x"1b1e",x"0756",x"051d",x"0820",x"19c2",x"1196",x"04af",x"1828",x"08ef",x"1198",x"1976",x"03f3",x"168e",x"1202",x"14c3",x"0a21",x"0b2a",x"0524",x"0080",x"1398",x"0432",x"1926",x"1f37",x"110c",x"127d",x"050f",x"001a",x"0797",x"16b8",x"1bdd",x"1710",x"0952",x"03ad",x"1ea1",x"10f6",x"1983",x"1e3a",x"0b66",x"1047",x"0839",x"0694",x"1970",x"05d8",x"0b42",x"1dfe",x"183c",x"020a",x"0233",x"1f62",x"1ed8",x"0500",x"1846",x"1b0d",x"0ae6",x"0419",x"045b",x"192f",x"0945",x"0ded",x"07fd",x"1669",x"1817",x"1fb3",x"09b6",x"0d18",x"05cd",x"1715",x"160d",x"0c42",x"0df8",x"0aa9",x"0a81",x"083a",x"0fed",x"0a34",x"0f80",x"0db9",x"077e",x"17fc",x"0a0e",x"1d64",x"1c87",
    --pkh
    x"79ba",x"7314",x"cebe",x"e997",x"f1ac",x"e68b",x"3987",x"187b", 
    x"7660",x"aa4b",x"974e",x"55f3",x"a7df",x"c8f0",x"00ca",x"c33a",
      --z
    x"f0b2",x"f504",x"5f43",x"c410",x"45cd",x"4811",x"7a44",x"9bfd", 
    x"b299",x"7709",x"e00d",x"3ad0",x"b7cd",x"6bbc",x"71e5",x"8c68",
    
    --SK--share1=======================================================================================================
--    --S polyvec 
--    x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
--    x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
--    x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
--    x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
--    x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
--    x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
--    x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
--    x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
    
--    x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
--    x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
--    x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
--    x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
--    x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
--    x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
--    x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
--    x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
    
--    x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
--    x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
--    x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
--    x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
--    x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
--    x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
--    x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
--    x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
    -- randmoly shared S polyvec
    
--    x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
--    x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
--    x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
    --rand shared
    x"00ae",x"0121",x"0833",x"0a79",x"132b",x"071f",x"0ecc",x"1e0b",x"12c1",x"0a64",x"1d2c",x"11f9",x"0c34",x"1cd6",x"0c61",x"1b51",x"0441",x"1532",x"1302",x"1d3b",x"098c",x"1acb",x"002b",x"190d",x"05be",x"1ed3",x"15f8",x"1f08",x"0ec8",x"0faa",x"1bab",x"02ba",x"1feb",x"1155",x"0ab6",x"0aa0",x"1206",x"0e9b",x"1aa9",x"1697",x"00ea",x"190d",x"0375",x"0b53",x"0fba",x"0920",x"0c61",x"1468",x"1b2e",x"02ba",x"1110",x"1625",x"06fe",x"155e",x"1256",x"0a96",x"0b99",x"1507",x"1954",x"17cc",x"141b",x"02a3",x"1e2f",x"164c",x"1831",x"1105",x"0ece",x"1655",x"1b17",x"12a3",x"1f7c",x"1548",x"0251",x"0889",x"1e17",x"066f",x"1cf1",x"1bcc",x"182a",x"1d3d",x"0a69",x"1014",x"1c47",x"0e69",x"00d4",x"02ac",x"1d11",x"0942",x"1bf0",x"12a0",x"06e6",x"12a8",x"1696",x"01a3",x"02c4",x"0d7d",x"166d",x"1d74",x"0f8e",x"12d5",x"18b7",x"0676",x"1540",x"1c24",x"0e8c",x"0152",x"1920",x"022a",x"0074",x"01b8",x"0151",x"1818",x"037c",x"1ad5",x"1d92",x"1e72",x"0b4c",x"04d9",x"17de",x"1899",x"06e4",x"198c",x"1bb0",x"17dc",x"0dfe",x"062c",x"06e0",x"03de",x"008a",x"0bfd",x"0260",x"1754",x"12a6",x"19fd",x"1e9f",x"0248",x"08ce",x"039b",x"0cd7",x"13ae",x"1ddb",x"1ecb",x"0429",x"1954",x"19a3",x"1883",x"0040",x"14d9",x"10dd",x"0a74",x"1730",x"0c64",x"0ae7",x"0703",x"1b0d",x"1fcb",x"0229",x"0141",x"02a7",x"1bb2",x"1960",x"1633",x"1689",x"1c77",x"0339",x"17d2",x"118c",x"0cab",x"0155",x"0224",x"08ec",x"1ef3",x"16fe",x"0e4d",x"1e19",x"174a",x"0b4e",x"1476",x"18e2",x"130a",x"19d8",x"1d58",x"050b",x"187a",x"1c67",x"1164",x"184f",x"0f47",x"19ef",x"1d82",x"06f8",x"16d4",x"0441",x"0f20",x"003f",x"0d1b",x"1082",x"0cee",x"1323",x"0e7b",x"03f8",x"133a",x"1a3e",x"0109",x"1256",x"1617",x"102f",x"0cb9",x"0859",x"14e9",x"1b28",x"094d",x"1287",x"056c",x"09d5",x"0cf8",x"0789",x"0330",x"1dcf",x"1d59",x"03ff",x"0de9",x"03e0",x"116c",x"016d",x"0cdc",x"0221",x"052b",x"0ba6",x"0622",x"09a3",x"00d5",x"0007",x"1c9c",x"0a2e",x"0f69",x"1a1e",x"0c60",x"014d",x"00ef",x"1606",x"13b3",x"11f8",x"1df5",x"1942",x"0938",x"0446",x"0ac7",x"15dc",x"1b58",x"042b",x"003f",x"1bde",x"1f2f",x"0e55",x"004d",x"13b9",x"137d",x"0458",x"0086",x"0fa4",x"1434",x"1959",x"1f2c",x"0cea",x"00ff",x"0f96",x"105e",x"1a84",x"043f",x"088e",x"15d6",x"155c",x"1013",x"0f93",x"1a26",x"0c2b",x"10d5",x"120a",x"1d3d",x"114b",x"1e3a",x"0ba3",x"07ff",x"0fea",x"072c",x"1ea6",x"06a4",x"06bb",x"086a",x"000f",x"0baf",x"06a1",x"130e",x"1940",x"0e0f",x"183d",x"1e9f",x"10e1",x"0a3a",x"0bcd",x"01c2",x"08f8",x"04e9",x"0bb7",x"1ab5",x"103b",x"10c4",x"1b09",x"1b99",x"10bb",x"1a0a",x"19e8",x"164f",x"14d8",x"057b",x"1059",x"0c7c",x"1d04",x"08ff",x"1443",x"18d7",x"0408",x"13f6",x"14f1",x"0348",x"01bc",x"1ff1",x"18f5",x"102b",x"1698",x"02d8",x"0b02",x"1e6a",x"148f",x"0564",x"1c88",x"1565",x"0b28",x"0424",x"1a66",x"0902",x"1482",x"0ba2",x"1587",x"084d",x"1e92",x"0561",x"0042",x"00c2",x"0a11",x"1c1d",x"13ab",x"04d2",x"0d77",x"01fc",x"1d9c",x"054a",x"0734",x"08c3",x"091a",x"1cc5",x"1a2e",x"1c47",x"082f",x"1aa8",x"17a8",x"0f9d",x"0b0e",x"10bf",x"1f33",x"06ac",x"03f9",x"1bab",x"08d4",x"0d07",x"0f31",x"13e0",x"0be1",x"12b4",x"1980",x"11fc",x"1e5a",x"1f09",x"1a42",x"1fc5",x"119b",x"041b",x"16e8",x"0c45",x"099d",x"1a95",x"0f1a",x"1251",x"1868",x"1ab0",x"130f",x"1391",x"0a01",x"0335",x"1565",x"1240",x"08ef",x"020d",x"1bb1",x"0113",x"0605",x"099d",x"1ffa",x"1268",x"1b0f",x"06d8",x"1dda",x"0092",x"15dc",x"1990",x"1999",x"1a3e",x"1320",x"10a9",x"1047",x"1307",x"12cf",x"0de2",x"1107",x"0920",x"0a26",x"12b7",x"0132",x"1928",x"1a5c",x"1861",x"0d1c",x"1b05",x"1450",x"1850",x"06c8",x"1d9b",x"1977",x"18ec",x"042b",x"03e5",x"1e5a",x"1820",x"0eff",x"1219",x"0950",x"0b2f",x"1d99",x"119a",x"0d9f",x"0bfd",x"07e7",x"0e4a",x"1390",x"1827",x"1742",x"1b02",x"0001",x"0e92",x"0e23",x"0d8d",x"1e47",x"0bbf",x"0195",x"1cae",x"06bb",x"0954",x"15b9",x"04c7",x"0657",x"199d",x"096d",x"13e0",x"132d",x"141d",x"07a9",x"1d9f",x"113f",x"0d81",x"0f28",x"1e93",x"08d1",x"048a",x"1dfc",x"17c1",x"1a5d",x"11c6",x"114e",x"1349",x"1e2d",x"00bd",x"08fb",x"0942",x"1231",x"1beb",x"0031",x"0faf",x"0cb2",x"06c7",x"0758",x"14de",x"0146",x"13e0",x"02ac",x"1e6b",x"1648",x"1dbc",x"0e37",x"0ea7",x"0335",x"0469",x"1702",x"06ba",x"1d41",x"124b",x"0df3",x"00af",x"018f",x"00d3",x"082b",x"1cbf",x"0723",x"1bf6",x"1dc9",x"0ca7",x"154a",x"061c",x"1406",x"0989",x"1cc9",x"0f46",x"12d0",x"06e9",x"025d",x"104d",x"00c4",x"1013",x"1a2c",x"10d7",x"1a81",x"0dbd",x"0edb",x"097d",x"022c",x"145a",x"0d23",x"04e0",x"0ba8",x"0355",x"0112",x"1208",x"0fea",x"0a1d",x"16bb",x"1dc8",x"1165",x"0e13",x"1f0e",x"031c",x"13c5",x"1b87",x"1765",x"1c41",x"171f",x"14d0",x"0ade",x"0465",x"0189",x"0638",x"0f19",x"0a36",x"1a30",x"1328",x"1cf8",x"104e",x"1adf",x"0758",x"1e58",x"00ee",x"1ae0",x"098f",x"1f88",x"1b03",x"09f7",x"01b4",x"09d2",x"1a7e",x"1d1e",x"0c29",x"0ec8",x"0abc",x"166e",x"0a80",x"166e",x"1e27",x"1193",x"042b",x"1fc8",x"141b",x"015a",x"1a74",x"1956",x"091a",x"14b1",x"065a",x"1f8a",x"0e69",x"1954",x"1f48",x"10ae",x"1c85",x"0542",x"1e7a",x"1893",x"1bea",x"04ed",x"17bb",x"06f8",x"1cdb",x"0391",x"0976",x"0b39",x"0ae7",x"0ddd",x"0a2d",x"15c3",x"175f",x"13ab",x"0239",x"0efe",x"09ef",x"1382",x"13a8",x"18c3",x"10c5",x"098c",x"13e9",x"0f84",x"1455",x"1d2f",x"0c71",x"1fd6",x"02c4",x"02ac",x"1205",x"0303",x"0e0c",x"091c",x"1e58",x"1a59",x"1333",x"1b3a",x"1e91",x"1ae7",x"12dd",x"0630",x"0f3c",x"0bf4",x"1fdc",x"0a98",x"0873",x"1c66",x"18ef",x"03ae",x"00c2",x"1286",x"186a",x"1a4e",x"0d87",x"0890",x"11f6",x"08d6",x"0658",x"1919",x"141a",x"07e5",x"028c",x"1d8b",x"1cd7",x"07c3",x"18f6",x"0437",x"1425",x"1b5e",x"0d82",x"04e2",x"18a8",x"1ae1",x"17df",x"063d",x"0e69",x"1b52",x"07d8",x"1712",x"0e67",x"068b",x"1c0e",x"0973",x"0dfe",x"0b3c",x"15df",x"14d7",x"1add",x"1f7f",x"0c69",x"1bcd",x"06dc",x"00ca",x"0ef6",x"0d83",x"1af2",x"1fe4",x"186a",x"0949",x"0423",x"08f1",x"16af",x"1c53",x"015d",x"0f0c",x"067e",x"01c6",x"149c",x"0fbc",x"17c6",x"196d",x"0690",x"1a28",x"14bf",x"0203",x"07c5",x"1df7",x"1dcd",x"00a0",x"0128",x"1aff",x"07bb",x"04f1",x"151c",x"1be8",x"1ba4",x"06d1",x"16bc",x"1213",x"1801",x"0996",x"07e8",x"004b",x"1648",x"12e7",x"1a31",x"08ed",x"09f3",x"13bd",x"1206",x"1557",x"157d",x"17c5",x"1014",x"15cb",x"107f",x"1248",x"1882",x"0803",x"15f0",x"029d",x"037b",
    --PKH
    x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
    x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
   
    --Z
    x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
    x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",

    --cipher = (Bp, cm)=========================================================
    --Bp
    -----Bp0
    x"5d4d", x"4b2b", x"29bf", x"93ef", x"4362", x"3017", x"470f", x"7c76", 
    x"a8a3", x"0a2a", x"1cf0", x"63cd", x"57f2", x"6440", x"ef29", x"ee31", 
    x"6b39", x"1367", x"0b76", x"84bb", x"05b4", x"a944", x"c640", x"1090", 
    x"11ad", x"07c6", x"320d", x"fac0", x"2a8d", x"60bc", x"0dc5", x"f351", 
    x"06e6", x"09c5", x"f254", x"cf60", x"0bbb", x"1dfd", x"d797", x"7543", 
    x"26e6", x"7eb8", x"9b05", x"fc42", x"bedf", x"08e2", x"a01e", x"7020", 
    x"633b", x"0dce", x"e876", x"05ca", x"1927", x"a0db", x"92db", x"feb4", 
    x"9059", x"baab", x"8562", x"1f7a", x"19aa", x"ff63", x"fa63", x"b212", 
    x"3f3f", x"1072", x"c5f2", x"802c", x"5029", x"4309", x"74d6", x"233f", 
    x"8731", x"e3d7", x"9c98", x"03f8", x"862f", x"f4d3", x"523b", x"f556", 
    x"50c2", x"c0ba", x"2708", x"5e45", x"54d8", x"ddf7", x"c705", x"1a5f", 
    x"b37c", x"573f", x"1f1c", x"e276", x"4c0d", x"12f9", x"0ce7", x"bde4", 
    x"754a", x"4894", x"ddea", x"1161", x"fe9b", x"0f27", x"3c8b", x"eba5", 
    x"4a80", x"8054", x"1ffc", x"e844", x"014b", x"6df2", x"ba76", x"6eb8", 
    x"75ff", x"aeeb", x"8a65", x"f5f2", x"8c8a", x"623e", x"f35a", x"b231", 
    x"3439", x"655f", x"63af", x"eb21", x"45cd", x"18dc", x"e07a", x"694e", 
    x"72ab", x"0288", x"1c6c", x"c6d0", x"3786", x"3391", x"62b6", x"7700", 
    x"5cc9", x"f859", x"849c", x"0351", x"5153", x"2d2c", x"dc32", x"c092", 
    x"1214", x"d456", x"e2b6", x"574c", x"c244", x"86bf", x"5766", x"52e5", 
    x"f509", x"067a", x"ce33", x"44c6", x"bd3e", x"910f", x"fea9", x"c454",
    ------Bp1
    x"1a43", x"979b", x"f4cf", x"e140", x"077d", x"b04f", x"e0b3", x"d6cb", 
    x"0447", x"50b4", x"178d", x"4b85", x"913a", x"70af", x"5b74", x"2c5f", 
    x"ab0a", x"5968", x"4219", x"dd0c", x"4850", x"d460", x"ae14", x"d975", 
    x"d21f", x"0e9d", x"839e", x"a924", x"e1d0", x"8b44", x"2ccb", x"1c7d", 
    x"1225", x"c76d", x"9425", x"d858", x"52f0", x"ca2a", x"b725", x"6a17", 
    x"b515", x"6638", x"fa63", x"5563", x"8189", x"8ced", x"7536", x"6be4", 
    x"1785", x"c827", x"5704", x"d157", x"3d25", x"1e2a", x"4718", x"4683", 
    x"6272", x"4649", x"0b4c", x"4de3", x"15a7", x"5d98", x"5376", x"b42c", 
    x"d4c7", x"a2b9", x"d6b3", x"08f8", x"546b", x"2870", x"7e99", x"eba8", 
    x"e47e", x"538b", x"b82e", x"50d9", x"e37b", x"04e8", x"d315", x"f0d8", 
    x"8b2b", x"34bf", x"56ee", x"39fa", x"1b9f", x"7e0e", x"2bd5", x"b700", 
    x"6bf6", x"1398", x"d0e4", x"31a3", x"8a98", x"1d73", x"1141", x"c095", 
    x"9711", x"520e", x"4d9e", x"ca35", x"1486", x"5036", x"82b6", x"050a", 
    x"d6a3", x"e606", x"1e72", x"0643", x"5927", x"0d64", x"4340", x"c927", 
    x"5b28", x"669f", x"95fd", x"6c8d", x"39ad", x"9b44", x"15f4", x"3621", 
    x"be44", x"25c5", x"6dd8", x"6152", x"d1f2", x"2bd1", x"b384", x"e72d", 
    x"a039", x"8df0", x"0f75", x"0ca2", x"f8d1", x"074a", x"0949", x"b20e", 
    x"9fa7", x"6295", x"d5f8", x"1ccd", x"48c6", x"3c11", x"981e", x"f6e9", 
    x"4326", x"de2d", x"c5c5", x"4b7b", x"ff17", x"71f7", x"e7d7", x"b954", 
    x"18b0", x"0b8f", x"70b8", x"280b", x"97cc", x"cb1d", x"b8aa", x"c0e4",
    ------Bp2
    x"f456", x"8c24", x"97ee", x"3018", x"7b35", x"3185", x"66d7", x"ebe2", 
    x"8d95", x"3349", x"ac78", x"1d24", x"1205", x"c80b", x"4e05", x"b767", 
    x"a450", x"16d8", x"7883", x"28d7", x"d61e", x"cb74", x"f416", x"a1f4", 
    x"5ab4", x"3c5d", x"9f04", x"eaf2", x"5b52", x"494a", x"5c1f", x"7c71", 
    x"4c11", x"4060", x"3677", x"cc31", x"2955", x"1054", x"2d23", x"5847", 
    x"748d", x"f65a", x"66f3", x"119a", x"eee9", x"c731", x"5ac5", x"1214", 
    x"5a30", x"283d", x"df7d", x"59f2", x"a71d", x"865a", x"8b0f", x"8926", 
    x"bd3b", x"8799", x"ed72", x"dbd7", x"1357", x"0bf4", x"4bd8", x"c65c", 
    x"fa1b", x"82c8", x"e4cf", x"0b5b", x"c3b8", x"1d6f", x"8251", x"df47", 
    x"6c72", x"9ba6", x"9bdc", x"7e5e", x"cc9c", x"7940", x"e397", x"72c0", 
    x"a787", x"da03", x"e7ec", x"708b", x"b422", x"5729", x"3eca", x"59ba", 
    x"cf19", x"6c8f", x"1e44", x"bcd0", x"4f57", x"75b4", x"77dc", x"1fe7", 
    x"693e", x"980b", x"14c6", x"5ffb", x"1549", x"ebbf", x"5f00", x"a3cb", 
    x"b6ba", x"e180", x"44c9", x"a495", x"d1b8", x"15ab", x"c400", x"6c87", 
    x"3219", x"782c", x"5eb8", x"3c69", x"9736", x"f36d", x"e34d", x"16f2", 
    x"0eec", x"a8d1", x"f3be", x"52fa", x"ac57", x"395f", x"0946", x"0634", 
    x"c4ee", x"aebf", x"757c", x"a21a", x"2521", x"3203", x"8f7b", x"0b0f", 
    x"278b", x"b7b3", x"193d", x"4a14", x"217c", x"28da", x"594d", x"8d67", 
    x"71cd", x"0615", x"435b", x"9f93", x"ddfd", x"1647", x"88e5", x"1059", 
    x"26c6", x"a330", x"501d", x"dc28", x"de04", x"b534", x"d7b8", x"c9ff",
    
    --cm
    x"0405", x"1812", x"b0fe", x"d0fd", x"234c", x"9051", x"20e6", x"f845", 
    x"ef72", x"212e", x"1ad5", x"eea4", x"ad8f", x"82d1", x"eee0", x"1d63", 
    x"5e13", x"5453", x"e907", x"fa0a", x"2432", x"92f6", x"e436", x"bfa3", 
    x"23ee", x"9f9a", x"1d50", x"d8a2", x"8507", x"fd07", x"ee21", x"52ce", 
    x"4f5e", x"e6b4", x"4046", x"d9f1", x"dd95", x"263c", x"6093", x"8b41", 
    x"88ff", x"92ee", x"6665", x"8d30", x"55fa", x"1dea", x"77b7", x"d231", 
    x"54eb", x"9bb2", x"7a8c", x"29c8", x"4a5e", x"e92f", x"c527", x"c00d", 
    x"ddbb", x"2da6", x"5ee8", x"c709", x"1c3a", x"62be", x"7e2d", x"0c19",
    --end chipertext
    
    others=>x"0000"
    );
    

end decaps_tv_shared_pkg;

package body decaps_tv_shared_pkg is
end package body;
